module tb();
reg a,b;

  //Write Code Here
initial begin
a = 1'b1;
b = 1'b0;
#10 a = 1'b1;
    b = 1'b1;
#10 a = 1'b0;
    b = 1'b1;
#10 a = 1'b0;
    b = 1'b0;
#10 a = 1'b1;
    b = 1'b0;
#10 $finish;
end
endmodule